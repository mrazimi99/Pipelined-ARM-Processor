module WBstage (input clk, rst, input[31: 0] pc_in, output[31: 0] pc);

  assign pc = pc_in;

endmodule // WBstage
