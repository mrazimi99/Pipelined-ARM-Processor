module ControlUnit (input[1: 0] mode, input[3: 0] op_code, input s, output aluCommand,
                    output mem_read, mem_write, wb_en, is_imm, branch, status_en);

endmodule // ControlUnit
