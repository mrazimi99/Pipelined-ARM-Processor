module ConditionCheck (input[3: 0] cond, input [31 :0] status,output result);

endmodule // ConditionCheck
